{AlgoIndexGtl: 4d} => '{VetoMask:01b}',
