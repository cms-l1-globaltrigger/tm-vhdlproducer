{AlgoIndexRop:d} => a_b_p({AlgoIndexGtl:d}),
