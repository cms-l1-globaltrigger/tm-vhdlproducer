{%- block bxComb_loop %}
  {%- for bx1, bx2 in module.muonBxCombinations %}
calc_muon_charge_correlations_bx_{{ bx1 }}_bx_{{ bx2 }}_i: entity work.muon_charge_correlations
    port map(mu_bx_{{ bx1 }}, mu_bx_{{ bx2 }},
        ls_charcorr_double_bx_{{ bx1 }}_bx_{{ bx2 }}, os_charcorr_double_bx_{{ bx1 }}_bx_{{ bx2 }},
        ls_charcorr_triple_bx_{{ bx1 }}_bx_{{ bx2 }}, os_charcorr_triple_bx_{{ bx1 }}_bx_{{ bx2 }},
        ls_charcorr_quad_bx_{{ bx1 }}_bx_{{ bx2 }}, os_charcorr_quad_bx_{{ bx1 }}_bx_{{ bx2 }});
--
  {%-endfor%}
{%- endblock bxComb_loop %}

