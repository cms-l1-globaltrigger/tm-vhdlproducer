    signal diff_{ObjectType}_wsc_eta_bx_{Bx} : diff_2dim_integer_array(0 to nr_{ObjectType}_objects-1, 0 to nr_{ObjectType}_objects-1) := (others => (others => 0));
    signal diff_{ObjectType}_wsc_phi_bx_{Bx} : diff_2dim_integer_array(0 to nr_{ObjectType}_objects-1, 0 to nr_{ObjectType}_objects-1) := (others => (others => 0));
