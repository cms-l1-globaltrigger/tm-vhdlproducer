    signal {ObjectType}_eta_bx_{Bx} : diff_inputs_array(0 to nr_{ObjectType}_objects-1) := (others => (others => '0'));
    signal {ObjectType}_eta_common_bx_{Bx} : diff_inputs_array(0 to nr_{ObjectType}_objects-1) := (others => (others => '0'));
    signal {ObjectType}_phi_bx_{Bx} : diff_inputs_array(0 to nr_{ObjectType}_objects-1) := (others => (others => '0'));
    signal {ObjectType}_phi_common_bx_{Bx} : diff_inputs_array(0 to nr_{ObjectType}_objects-1) := (others => (others => '0'));
