-- future delta r condition
