{ConditionName}_i: muon_conditions
    generic map(nr_muon_objects, {NrTemplates:d}, {DoubleWsc}, {PtGeMode}, d_s_i_muon,
        (X"{PtThresholds[0]:04X}", X"{PtThresholds[1]:04X}", X"{PtThresholds[2]:04X}", X"{PtThresholds[3]:04X}"),
        ({EtaFullRange[0]}, {EtaFullRange[1]}, {EtaFullRange[2]}, {EtaFullRange[3]}),
        (X"{EtaW1UpperLimits[0]:04X}", X"{EtaW1UpperLimits[1]:04X}", X"{EtaW1UpperLimits[2]:04X}", X"{EtaW1UpperLimits[3]:04X}"), (X"{EtaW1LowerLimits[0]:04X}", X"{EtaW1LowerLimits[1]:04X}", X"{EtaW1LowerLimits[2]:04X}", X"{EtaW1LowerLimits[3]:04X}"),
        ({EtaW2Ignore[0]}, {EtaW2Ignore[1]}, {EtaW2Ignore[2]}, {EtaW2Ignore[3]}),
        (X"{EtaW2UpperLimits[0]:04X}", X"{EtaW2UpperLimits[1]:04X}", X"{EtaW2UpperLimits[2]:04X}", X"{EtaW2UpperLimits[3]:04X}"), (X"{EtaW2LowerLimits[0]:04X}", X"{EtaW2LowerLimits[1]:04X}", X"{EtaW2LowerLimits[2]:04X}", X"{EtaW2LowerLimits[3]:04X}"),
        ({PhiFullRange[0]}, {PhiFullRange[1]}, {PhiFullRange[2]}, {PhiFullRange[3]}),
        (X"{PhiW1UpperLimits[0]:04X}", X"{PhiW1UpperLimits[1]:04X}", X"{PhiW1UpperLimits[2]:04X}", X"{PhiW1UpperLimits[3]:04X}"), (X"{PhiW1LowerLimits[0]:04X}", X"{PhiW1LowerLimits[1]:04X}", X"{PhiW1LowerLimits[2]:04X}", X"{PhiW1LowerLimits[3]:04X}"),
        ({PhiW2Ignore[0]}, {PhiW2Ignore[1]}, {PhiW2Ignore[2]}, {PhiW2Ignore[3]}),
        (X"{PhiW2UpperLimits[0]:04X}", X"{PhiW2UpperLimits[1]:04X}", X"{PhiW2UpperLimits[2]:04X}", X"{PhiW2UpperLimits[3]:04X}"), (X"{PhiW2LowerLimits[0]:04X}", X"{PhiW2LowerLimits[1]:04X}", X"{PhiW2LowerLimits[2]:04X}", X"{PhiW2LowerLimits[3]:04X}"),
        ("{RequestedCharges[0]}", "{RequestedCharges[1]}", "{RequestedCharges[2]}", "{RequestedCharges[3]}"),
        (X"{QualityLuts[0]:04X}", X"{QualityLuts[1]:04X}", X"{QualityLuts[2]:04X}", X"{QualityLuts[3]:04X}"),
        (X"{IsolationLuts[0]:01X}", X"{IsolationLuts[1]:01X}", X"{IsolationLuts[2]:01X}", X"{IsolationLuts[3]:01X}"),
        "{RequestedChargeCorrelation}",
        {DiffEtaUpperLimit:d}, {DiffEtaLowerLimit:d}, {DiffPhiUpperLimit:d}, {DiffPhiLowerLimit:d})
    port map(lhc_clk, muon_bx_{Bx},
        ls_charcorr_double_bx_{Bx}, os_charcorr_double_bx_{Bx},
        ls_charcorr_triple_bx_{Bx}, os_charcorr_triple_bx_{Bx},
        ls_charcorr_quad_bx_{Bx}, os_charcorr_quad_bx_{Bx},
        diff_muon_wsc_eta_bx_{Bx}, diff_muon_wsc_phi_bx_{Bx},
        {ConditionName});
