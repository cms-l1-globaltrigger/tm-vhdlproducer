{AlgoIndexGtl: 4d} => '{FinorMask:01b}',
