    signal diff_{ObjectType1}_{ObjectType2}_eta_bx_{Bx1}_bx_{Bx2} : diff_2dim_integer_array(0 to nr_{ObjectType1}_objects-1, 0 to nr_{ObjectType2}_objects-1) := (others => (others => 0));
    signal diff_{ObjectType1}_{ObjectType2}_phi_bx_{Bx1}_bx_{Bx2} : diff_2dim_integer_array(0 to nr_{ObjectType1}_objects-1, 0 to nr_{ObjectType2}_objects-1) := (others => (others => 0));
