{AlgoIndexGtl: 4d} => X"{FinorVetoMasks:08X}",
