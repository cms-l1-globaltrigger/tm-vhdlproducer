    signal {AlgoName} : std_logic;
