{%- block signal_correlation_conditions_pt_eta_phi_cos_sin_loop %}
  {%- for o in module.correlationObjects %}
    {%- if o.is_calo_type %}
    signal {{ o.type|lower }}_pt_vector_bx_{{ o.bx }}: diff_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => (others => '0'));
    signal {{ o.type|lower }}_eta_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_phi_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_cos_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_sin_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal conv_{{ o.type|lower }}_cos_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal conv_{{ o.type|lower }}_sin_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_eta_conv_2_muon_eta_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_phi_conv_2_muon_phi_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    {%- elif o.is_muon_type %}
    signal {{ o.type|lower }}_pt_vector_bx_{{ o.bx }}: diff_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => (others => '0'));
    signal {{ o.type|lower }}_upt_vector_bx_{{ o.bx }}: diff_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => (others => '0'));
    signal {{ o.type|lower }}_eta_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_phi_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_cos_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_sin_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    {%- elif o.is_esums_type %}
    signal {{ o.type|lower }}_pt_vector_bx_{{ o.bx }}: diff_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => (others => '0'));
    signal {{ o.type|lower }}_phi_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_cos_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_sin_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal conv_{{ o.type|lower }}_cos_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal conv_{{ o.type|lower }}_sin_phi_bx_{{ o.bx }}: sin_cos_integer_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    signal {{ o.type|lower }}_phi_conv_2_muon_phi_integer_bx_{{ o.bx }}: diff_integer_inputs_array(0 to NR_{{ o.type|upper }}_OBJECTS-1) := (others => 0);
    {%- endif %}
  {%- endfor %}
{%- endblock signal_correlation_conditions_pt_eta_phi_cos_sin_loop %}
{# eof #}
