    signal {ConditionName} : std_logic;
