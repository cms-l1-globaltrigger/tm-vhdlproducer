{AlgoIndexRop:d} => a_a_f({AlgoIndexGtl:d}),
