{AlgoIndexRop:d} => a_a_p({AlgoIndexGtl:d}),
