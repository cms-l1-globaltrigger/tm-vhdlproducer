{AlgoIndexGtl: 4d} => X"{PrescaleFactor:08X}",
