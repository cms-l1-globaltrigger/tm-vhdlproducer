{AlgoName} <= {AlgoEquation};
algo({AlgoIndex:d}) <= {AlgoName};
