    signal pos_charge_single_bx_{Bx} : muon_charge_1_array;
    signal neg_charge_single_bx_{Bx} : muon_charge_1_array;
    signal eq_charge_double_bx_{Bx} : muon_charge_2_array;
    signal neq_charge_double_bx_{Bx} : muon_charge_2_array;
    signal eq_charge_triple_bx_{Bx} : muon_charge_3_array;
    signal neq_charge_triple_bx_{Bx} : muon_charge_3_array;
    signal eq_charge_quad_bx_{Bx} : muon_charge_4_array;
    signal pair_charge_quad_bx_{Bx} : muon_charge_4_array;
