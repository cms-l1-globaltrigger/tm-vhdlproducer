muon_charge_correlations_bx_{Bx}_i: muon_charge_correlations
    port map(muon_bx_{Bx},
        ls_charcorr_double_bx_{Bx}, os_charcorr_double_bx_{Bx},
        ls_charcorr_triple_bx_{Bx}, os_charcorr_triple_bx_{Bx},
        ls_charcorr_quad_bx_{Bx}, os_charcorr_quad_bx_{Bx});
