    signal ls_charcorr_double_bx_{Bx}, os_charcorr_double_bx_{Bx} : muon_charcorr_double_array;
    signal ls_charcorr_triple_bx_{Bx}, os_charcorr_triple_bx_{Bx} : muon_charcorr_triple_array;
    signal ls_charcorr_quad_bx_{Bx}, os_charcorr_quad_bx_{Bx} : muon_charcorr_quad_array;
