muon_charges_bx_{Bx}_i: muon_charges
    port map(muon_bx_{Bx}, pos_charge_single_bx_{Bx}, neg_charge_single_bx_{Bx},
        eq_charge_double_bx_{Bx}, neq_charge_double_bx_{Bx},
        eq_charge_triple_bx_{Bx}, neq_charge_triple_bx_{Bx},
        eq_charge_quad_bx_{Bx}, pair_charge_quad_bx_{Bx});
